LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- declaracao de entidade
ENTITY MEUCIRCUITO IS
	PORT (A, B, C: IN STD_LOGIC;
		X,Y: OUT STD_LOGIC;)
END MEUCIRCUITO;

-- circuito 1

ARCHITECTURE MEUCIRCUITO_ARCH OF MEUCIRCUITO IS
BEGIN 
	X <= (NOT(A) AND C) OR (A AND B);
	Y <= (NOT(A) AND C) OR (A AND B);
END MEUCIRCUITO_ARCH;

-- circuito 2

ARCHITECTURE MEUCIRCUITO_ARCH2 OF MEUCIRCUITO IS
SIGNAL FIO1, FIO2: STD_LOGIC;
BEGIN
	FIO1 <= NOT(A) AND C;
	FIO2 <= A AND B;
	X <= FIO1 OR FIO2;
	Y <= FIO1 OR NOT(FIO2);
END MEUCIRCUITO_ARCH2;
