LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY HELLOWORLD IS
	PORT(A, B, Cin: IN STD_LOGIC;
	     S, Cout: OUT STD_LOGIC);
END HELLOWORLD;

ARCHITECTURE HELLOWORLD_EXE OF HELLOWORLD IS
BEGIN
	S <= A XOR B XOR Cin;
	Cout <= (A AND B) OR (A AND Cin) OR (B AND Cin);
END HELLOWORLD_EXE;


	 